module DMUXzm16z_workaround (clk, rst, Selector, Disable, Output_1, Output_2, Output_3, Output_4, Output_5, Output_6, Output_7, Output_8, Output_9, Output_10, Output_11, Output_12, Output_13, Output_14, Output_15, Output_16);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] Selector;
  input  wire [0:0] Disable;
  output  wire [0:0] Output_1;
  output  wire [0:0] Output_2;
  output  wire [0:0] Output_3;
  output  wire [0:0] Output_4;
  output  wire [0:0] Output_5;
  output  wire [0:0] Output_6;
  output  wire [0:0] Output_7;
  output  wire [0:0] Output_8;
  output  wire [0:0] Output_9;
  output  wire [0:0] Output_10;
  output  wire [0:0] Output_11;
  output  wire [0:0] Output_12;
  output  wire [0:0] Output_13;
  output  wire [0:0] Output_14;
  output  wire [0:0] Output_15;
  output  wire [0:0] Output_16;

  TC_Splitter8 # (.UUID(64'd2501185698665852659 ^ UUID)) Splitter8_0 (.in(wire_14), .out0(wire_0), .out1(wire_15), .out2(wire_9), .out3(wire_2), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd3051034902902567548 ^ UUID)) Decoder3_1 (.dis(wire_24), .sel0(wire_0), .sel1(wire_15), .sel2(wire_9), .out0(wire_19), .out1(wire_5), .out2(wire_20), .out3(wire_6), .out4(wire_10), .out5(wire_18), .out6(wire_11), .out7(wire_13));
  TC_Decoder3 # (.UUID(64'd3176597986420345467 ^ UUID)) Decoder3_2 (.dis(wire_23), .sel0(wire_0), .sel1(wire_15), .sel2(wire_9), .out0(wire_4), .out1(wire_16), .out2(wire_21), .out3(wire_17), .out4(wire_8), .out5(wire_1), .out6(wire_12), .out7(wire_3));
  TC_Not # (.UUID(64'd3649176789582710296 ^ UUID), .BIT_WIDTH(64'd1)) Not_3 (.in(wire_2), .out(wire_22));
  TC_Switch # (.UUID(64'd2627742891582984678 ^ UUID), .BIT_WIDTH(64'd1)) Output1z_4 (.en(wire_3), .in(wire_3), .out(Output_9));
  TC_Switch # (.UUID(64'd2959290984966874439 ^ UUID), .BIT_WIDTH(64'd1)) Output1z_5 (.en(wire_12), .in(wire_12), .out(Output_10));
  TC_Switch # (.UUID(64'd3287414910794005956 ^ UUID), .BIT_WIDTH(64'd1)) Output1z_6 (.en(wire_1), .in(wire_1), .out(Output_11));
  TC_Switch # (.UUID(64'd1180559238184509638 ^ UUID), .BIT_WIDTH(64'd1)) Output1z_7 (.en(wire_8), .in(wire_8), .out(Output_12));
  TC_Switch # (.UUID(64'd3756066530922898251 ^ UUID), .BIT_WIDTH(64'd1)) Output1z_8 (.en(wire_17), .in(wire_17), .out(Output_13));
  TC_Switch # (.UUID(64'd845184652869544769 ^ UUID), .BIT_WIDTH(64'd1)) Output1z_9 (.en(wire_21), .in(wire_21), .out(Output_14));
  TC_Switch # (.UUID(64'd816809522013653411 ^ UUID), .BIT_WIDTH(64'd1)) Output1z_10 (.en(wire_16), .in(wire_16), .out(Output_15));
  TC_Switch # (.UUID(64'd2821416941940642917 ^ UUID), .BIT_WIDTH(64'd1)) Output1z_11 (.en(wire_4), .in(wire_4), .out(Output_16));
  TC_Switch # (.UUID(64'd4353151609242476992 ^ UUID), .BIT_WIDTH(64'd1)) Output1z_12 (.en(wire_13), .in(wire_13), .out(Output_1));
  TC_Switch # (.UUID(64'd2291511641141839562 ^ UUID), .BIT_WIDTH(64'd1)) Output1z_13 (.en(wire_11), .in(wire_11), .out(Output_2));
  TC_Switch # (.UUID(64'd997920623655650288 ^ UUID), .BIT_WIDTH(64'd1)) Output1z_14 (.en(wire_18), .in(wire_18), .out(Output_3));
  TC_Switch # (.UUID(64'd1149460066355519615 ^ UUID), .BIT_WIDTH(64'd1)) Output1z_15 (.en(wire_10), .in(wire_10), .out(Output_4));
  TC_Switch # (.UUID(64'd4212664422248886661 ^ UUID), .BIT_WIDTH(64'd1)) Output1z_16 (.en(wire_6), .in(wire_6), .out(Output_5));
  TC_Switch # (.UUID(64'd3579460137179712060 ^ UUID), .BIT_WIDTH(64'd1)) Output1z_17 (.en(wire_20), .in(wire_20), .out(Output_6));
  TC_Switch # (.UUID(64'd4210674212345144653 ^ UUID), .BIT_WIDTH(64'd1)) Output1z_18 (.en(wire_5), .in(wire_5), .out(Output_7));
  TC_Switch # (.UUID(64'd3072089910523482094 ^ UUID), .BIT_WIDTH(64'd1)) Output1z_19 (.en(wire_19), .in(wire_19), .out(Output_8));
  OR # (.UUID(64'd2893939579020398837 ^ UUID)) OR_20 (.clk(clk), .rst(rst), .Input_1(wire_2), .Input_2(wire_7), .Output(wire_24));
  OR # (.UUID(64'd2274188548802102818 ^ UUID)) OR_21 (.clk(clk), .rst(rst), .Input_1(wire_22), .Input_2(wire_7), .Output(wire_23));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  assign wire_7 = Disable;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [7:0] wire_14;
  assign wire_14 = Selector;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;

endmodule
