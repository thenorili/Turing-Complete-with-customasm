module MUXzm16zp (clk, rst, \0 , \1 , \2 , \3 , \4 , \5 , \6 , \7 , Selector, \15 , \14 , \13 , \12 , \11 , \10 , \9 , \8 , Disable, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] \0 ;
  input  wire [7:0] \1 ;
  input  wire [7:0] \2 ;
  input  wire [7:0] \3 ;
  input  wire [7:0] \4 ;
  input  wire [7:0] \5 ;
  input  wire [7:0] \6 ;
  input  wire [7:0] \7 ;
  input  wire [7:0] Selector;
  input  wire [7:0] \15 ;
  input  wire [7:0] \14 ;
  input  wire [7:0] \13 ;
  input  wire [7:0] \12 ;
  input  wire [7:0] \11 ;
  input  wire [7:0] \10 ;
  input  wire [7:0] \9 ;
  input  wire [7:0] \8 ;
  input  wire [0:0] Disable;
  output  wire [7:0] Output;

  TC_Switch # (.UUID(64'd3191703730251323901 ^ UUID), .BIT_WIDTH(64'd8)) Output8z_0 (.en(wire_6), .in(wire_0), .out(Output));
  TC_Splitter8 # (.UUID(64'd4005357342071797364 ^ UUID)) Splitter8_1 (.in(wire_12), .out0(), .out1(), .out2(), .out3(wire_4), .out4(), .out5(), .out6(), .out7());
  TC_Not # (.UUID(64'd4348972499109896650 ^ UUID), .BIT_WIDTH(64'd1)) Not_2 (.in(wire_4), .out(wire_3));
  TC_Not # (.UUID(64'd519778269274372978 ^ UUID), .BIT_WIDTH(64'd1)) Not_3 (.in(wire_7), .out(wire_6));
  MUXzm8zp # (.UUID(64'd3055454744049391241 ^ UUID)) MUXzm8zp_4 (.clk(clk), .rst(rst), .\0 (wire_17), .\1 (wire_22), .\2 (wire_21), .\3 (wire_15), .\4 (wire_2), .\5 (wire_9), .\6 (wire_18), .\7 (wire_11), .Selector(wire_12), .Disable(wire_23), .Output(wire_0_1));
  MUXzm8zp # (.UUID(64'd3482936192979053147 ^ UUID)) MUXzm8zp_5 (.clk(clk), .rst(rst), .\0 (wire_20), .\1 (wire_13), .\2 (wire_14), .\3 (wire_5), .\4 (wire_8), .\5 (wire_16), .\6 (wire_19), .\7 (wire_1), .Selector(wire_12), .Disable(wire_10), .Output(wire_0_0));
  OR # (.UUID(64'd1515119195311848162 ^ UUID)) OR_6 (.clk(clk), .rst(rst), .Input_1(wire_4), .Input_2(wire_7), .Output(wire_23));
  OR # (.UUID(64'd1103179269122331715 ^ UUID)) OR_7 (.clk(clk), .rst(rst), .Input_1(wire_7), .Input_2(wire_3), .Output(wire_10));

  wire [7:0] wire_0;
  wire [7:0] wire_0_0;
  wire [7:0] wire_0_1;
  assign wire_0 = wire_0_0|wire_0_1;
  wire [7:0] wire_1;
  assign wire_1 = \15 ;
  wire [7:0] wire_2;
  assign wire_2 = \4 ;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [7:0] wire_5;
  assign wire_5 = \11 ;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  assign wire_7 = Disable;
  wire [7:0] wire_8;
  assign wire_8 = \12 ;
  wire [7:0] wire_9;
  assign wire_9 = \5 ;
  wire [0:0] wire_10;
  wire [7:0] wire_11;
  assign wire_11 = \7 ;
  wire [7:0] wire_12;
  assign wire_12 = Selector;
  wire [7:0] wire_13;
  assign wire_13 = \9 ;
  wire [7:0] wire_14;
  assign wire_14 = \10 ;
  wire [7:0] wire_15;
  assign wire_15 = \3 ;
  wire [7:0] wire_16;
  assign wire_16 = \13 ;
  wire [7:0] wire_17;
  assign wire_17 = \0 ;
  wire [7:0] wire_18;
  assign wire_18 = \6 ;
  wire [7:0] wire_19;
  assign wire_19 = \14 ;
  wire [7:0] wire_20;
  assign wire_20 = \8 ;
  wire [7:0] wire_21;
  assign wire_21 = \2 ;
  wire [7:0] wire_22;
  assign wire_22 = \1 ;
  wire [0:0] wire_23;

endmodule
