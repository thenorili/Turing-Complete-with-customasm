module LEGz_06z_callret (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_IOSwitch # (.UUID(64'd4389593845 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_0 (.in(wire_0), .en(wire_40), .out(arch_output_value));
  TC_Switch # (.UUID(64'd438959385 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_1 (.en(wire_62), .in(arch_input_value), .out(wire_5));
  TC_Counter # (.UUID(64'd4227818422159936411 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd4)) Counter8_2 (.clk(clk), .rst(rst), .save(wire_64), .in(wire_0), .out(wire_74));
  TC_Register # (.UUID(64'd4607782328979482347 ^ UUID), .BIT_WIDTH(64'd8)) Register8_3 (.clk(clk), .rst(rst), .load(wire_18), .save(wire_47), .in(wire_0), .out(wire_35));
  TC_Register # (.UUID(64'd2654441428106189356 ^ UUID), .BIT_WIDTH(64'd8)) Register8_4 (.clk(clk), .rst(rst), .load(wire_53), .save(wire_37), .in(wire_0), .out(wire_31));
  TC_Register # (.UUID(64'd1441950349091143385 ^ UUID), .BIT_WIDTH(64'd8)) Register8_5 (.clk(clk), .rst(rst), .load(wire_50), .save(wire_33), .in(wire_0), .out(wire_56));
  TC_Register # (.UUID(64'd3728739506887436998 ^ UUID), .BIT_WIDTH(64'd8)) Register8_6 (.clk(clk), .rst(rst), .load(wire_36), .save(wire_60), .in(wire_0), .out(wire_9));
  TC_Register # (.UUID(64'd813762756125550530 ^ UUID), .BIT_WIDTH(64'd8)) Register8_7 (.clk(clk), .rst(rst), .load(wire_32), .save(wire_2), .in(wire_0), .out(wire_1));
  TC_Register # (.UUID(64'd4029391467152470696 ^ UUID), .BIT_WIDTH(64'd8)) Register8_8 (.clk(clk), .rst(rst), .load(wire_48), .save(wire_42), .in(wire_0), .out(wire_55));
  TC_Decoder3 # (.UUID(64'd3632482315835268131 ^ UUID)) Decoder3_9 (.dis(wire_72), .sel0(wire_71), .sel1(wire_73), .sel2(wire_38), .out0(wire_47), .out1(wire_37), .out2(wire_33), .out3(wire_60), .out4(wire_2), .out5(wire_42), .out6(wire_63), .out7(wire_21));
  TC_Splitter8 # (.UUID(64'd2588566827510959189 ^ UUID)) Splitter8_10 (.in(wire_25[7:0]), .out0(wire_71), .out1(wire_73), .out2(wire_38), .out3(wire_34), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd850112712224890741 ^ UUID)) Splitter8_11 (.in(wire_14[7:0]), .out0(), .out1(), .out2(), .out3(), .out4(), .out5(wire_4), .out6(wire_23), .out7(wire_11));
  TC_Mux # (.UUID(64'd2967387940270423087 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_12 (.sel(wire_11), .in0(wire_69), .in1(wire_16[7:0]), .out(wire_15));
  TC_Mux # (.UUID(64'd4133036621474758973 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_13 (.sel(wire_23), .in0(wire_10), .in1(wire_6[7:0]), .out(wire_13));
  TC_Mux # (.UUID(64'd4189709243187177903 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_14 (.sel(wire_4), .in0(wire_44), .in1(wire_25[7:0]), .out(wire_0));
  TC_Decoder3 # (.UUID(64'd4528304914669755354 ^ UUID)) Decoder3_15 (.dis(wire_67), .sel0(wire_71), .sel1(wire_73), .sel2(wire_38), .out0(wire_26), .out1(wire_29), .out2(wire_65), .out3(wire_27), .out4(wire_17), .out5(wire_24), .out6(wire_30), .out7(wire_40));
  TC_Not # (.UUID(64'd676189359525278885 ^ UUID), .BIT_WIDTH(64'd1)) Not_16 (.in(wire_34), .out(wire_68));
  TC_Ram # (.UUID(64'd4372783762123074173 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd256)) Ram_17 (.clk(clk), .rst(rst), .load(wire_49), .save(wire_24), .address({{24{1'b0}}, wire_45 }), .in0({{56{1'b0}}, wire_0 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_3), .out1(), .out2(), .out3());
  TC_Register # (.UUID(64'd3855708699894118692 ^ UUID), .BIT_WIDTH(64'd8)) Register8_18 (.clk(clk), .rst(rst), .load(wire_52), .save(wire_21), .in(wire_0), .out(wire_66));
  TC_Register # (.UUID(64'd2875837445672808175 ^ UUID), .BIT_WIDTH(64'd8)) Register8_19 (.clk(clk), .rst(rst), .load(wire_8), .save(wire_26), .in(wire_0), .out(wire_7));
  TC_Register # (.UUID(64'd2275915933328980784 ^ UUID), .BIT_WIDTH(64'd8)) Register8_20 (.clk(clk), .rst(rst), .load(wire_28), .save(wire_29), .in(wire_0), .out(wire_43));
  TC_Register # (.UUID(64'd2198714164874018182 ^ UUID), .BIT_WIDTH(64'd8)) Register8_21 (.clk(clk), .rst(rst), .load(wire_57), .save(wire_17), .in(wire_0), .out(wire_45));
  TC_Register # (.UUID(64'd1456120796309230852 ^ UUID), .BIT_WIDTH(64'd8)) Register8_22 (.clk(clk), .rst(rst), .load(wire_59), .save(wire_63), .in(wire_0), .out(wire_39));
  TC_Constant # (.UUID(64'd897712722238026467 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_23 (.out(wire_57));
  TC_Switch # (.UUID(64'd35036273375025196 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_24 (.en(wire_46), .in(wire_45), .out(wire_19));
  TC_Program # (.UUID(64'd2945955032425777044 ^ UUID), .WORD_WIDTH(64'd8), .DEFAULT_FILE_NAME("Program_28E2227E60034794.w8.bin"), .ARG_SIG("Program_28E2227E60034794=%s")) Program_25 (.clk(clk), .rst(rst), .address({{8{1'b0}}, wire_74 }), .out0(wire_14), .out1(wire_16), .out2(wire_6), .out3(wire_25));
  TC_Register # (.UUID(64'd467538734190536617 ^ UUID), .BIT_WIDTH(64'd8)) Register8_26 (.clk(clk), .rst(rst), .load(wire_54), .save(wire_27), .in(wire_0), .out(wire_61));
  TC_Register # (.UUID(64'd1607121337331166466 ^ UUID), .BIT_WIDTH(64'd8)) Register8_27 (.clk(clk), .rst(rst), .load(wire_51), .save(wire_30), .in(wire_0), .out(wire_22));
  CONDzmLEG # (.UUID(64'd3310312642247156829 ^ UUID)) CONDzmLEG_28 (.clk(clk), .rst(rst), .Input_1(wire_15), .Input_2(wire_13), .Opcode(wire_14[7:0]), .Output(wire_58));
  ALUzmLEGzm16 # (.UUID(64'd3486083726480225081 ^ UUID)) ALUzmLEGzm16_29 (.clk(clk), .rst(rst), .Input_1(wire_15), .Input_2(wire_13), .Opcode(wire_14[7:0]), .Output(wire_44));
  OR # (.UUID(64'd1225838809174928741 ^ UUID)) OR_30 (.clk(clk), .rst(rst), .Input_1(wire_4), .Input_2(wire_34), .Output(wire_72));
  OR # (.UUID(64'd2082960413066559696 ^ UUID)) OR_31 (.clk(clk), .rst(rst), .Input_1(wire_68), .Input_2(wire_4), .Output(wire_67));
  MUXzm16zp # (.UUID(64'd319829999529271899 ^ UUID)) MUXzm16zp_32 (.clk(clk), .rst(rst), .\0 (wire_35), .\1 (wire_31), .\2 (wire_56), .\3 (wire_9), .\4 (wire_1), .\5 (wire_55), .\6 (wire_39), .\7 (wire_66), .Selector(wire_16[7:0]), .\15 (wire_5), .\14 (wire_22), .\13 (wire_3[7:0]), .\12 (wire_19), .\11 (wire_61), .\10 ({{7{1'b0}}, wire_12 }), .\9 (wire_43), .\8 (wire_7), .Disable(1'd0), .Output(wire_69));
  MUXzm16zp # (.UUID(64'd2651032360632107951 ^ UUID)) MUXzm16zp_33 (.clk(clk), .rst(rst), .\0 (wire_35), .\1 (wire_31), .\2 (wire_56), .\3 (wire_9), .\4 (wire_1), .\5 (wire_55), .\6 (wire_39), .\7 (wire_66), .Selector(wire_6[7:0]), .\15 (wire_5), .\14 (wire_22), .\13 (wire_3[7:0]), .\12 (wire_19), .\11 (wire_61), .\10 ({{7{1'b0}}, wire_12 }), .\9 (wire_43), .\8 (wire_7), .Disable(1'd0), .Output(wire_10));
  DMUXzm16z_workaround # (.UUID(64'd3328331167516938516 ^ UUID)) DMUXzm16z_workaround_34 (.clk(clk), .rst(rst), .Selector(wire_6[7:0]), .Disable(1'd0), .Output_1(wire_52_0), .Output_2(wire_59_1), .Output_3(wire_48_0), .Output_4(wire_32_0), .Output_5(wire_36_0), .Output_6(wire_50_0), .Output_7(wire_53_0), .Output_8(wire_18_1), .Output_9(wire_62_0), .Output_10(wire_51_0), .Output_11(wire_49_0), .Output_12(wire_46_0), .Output_13(wire_54_0), .Output_14(wire_70_1), .Output_15(wire_28_0), .Output_16(wire_8_0));
  DMUXzm16z_workaround # (.UUID(64'd1462152971226604546 ^ UUID)) DMUXzm16z_workaround_35 (.clk(clk), .rst(rst), .Selector(wire_16[7:0]), .Disable(1'd0), .Output_1(wire_52_1), .Output_2(wire_59_0), .Output_3(wire_48_1), .Output_4(wire_32_1), .Output_5(wire_36_1), .Output_6(wire_50_1), .Output_7(wire_53_1), .Output_8(wire_18_0), .Output_9(wire_62_1), .Output_10(wire_51_1), .Output_11(wire_49_1), .Output_12(wire_46_1), .Output_13(wire_54_1), .Output_14(wire_70_0), .Output_15(wire_28_1), .Output_16(wire_8_1));
  AND # (.UUID(64'd2224082151904094725 ^ UUID)) AND_36 (.clk(clk), .rst(rst), .Input_1(wire_4), .Input_2(wire_58), .Output(wire_20));
  TC_Halt # (.UUID(64'd4342208852562261490 ^ UUID)) Halt_37 (.clk(clk), .rst(rst), .en(wire_41));
  TC_Switch # (.UUID(64'd2126690747936412766 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_38 (.en(wire_40), .in(wire_40), .out(wire_41));
  OR # (.UUID(64'd4425575856016504479 ^ UUID)) OR_39 (.clk(clk), .rst(rst), .Input_1(wire_20), .Input_2(wire_65), .Output(wire_64));

  wire [7:0] wire_0;
  wire [7:0] wire_1;
  wire [0:0] wire_2;
  wire [63:0] wire_3;
  wire [0:0] wire_4;
  wire [7:0] wire_5;
  wire [63:0] wire_6;
  wire [7:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_8_0;
  wire [0:0] wire_8_1;
  assign wire_8 = wire_8_0|wire_8_1;
  wire [7:0] wire_9;
  wire [7:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  assign wire_12 = 0;
  wire [7:0] wire_13;
  wire [63:0] wire_14;
  wire [7:0] wire_15;
  wire [63:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_18_0;
  wire [0:0] wire_18_1;
  assign wire_18 = wire_18_0|wire_18_1;
  wire [7:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [7:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [63:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_28_0;
  wire [0:0] wire_28_1;
  assign wire_28 = wire_28_0|wire_28_1;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [7:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_32_0;
  wire [0:0] wire_32_1;
  assign wire_32 = wire_32_0|wire_32_1;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [7:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_36_0;
  wire [0:0] wire_36_1;
  assign wire_36 = wire_36_0|wire_36_1;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [7:0] wire_39;
  wire [0:0] wire_40;
  assign arch_output_enable = wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [7:0] wire_43;
  wire [7:0] wire_44;
  wire [7:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_46_0;
  wire [0:0] wire_46_1;
  assign wire_46 = wire_46_0|wire_46_1;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_48_0;
  wire [0:0] wire_48_1;
  assign wire_48 = wire_48_0|wire_48_1;
  wire [0:0] wire_49;
  wire [0:0] wire_49_0;
  wire [0:0] wire_49_1;
  assign wire_49 = wire_49_0|wire_49_1;
  wire [0:0] wire_50;
  wire [0:0] wire_50_0;
  wire [0:0] wire_50_1;
  assign wire_50 = wire_50_0|wire_50_1;
  wire [0:0] wire_51;
  wire [0:0] wire_51_0;
  wire [0:0] wire_51_1;
  assign wire_51 = wire_51_0|wire_51_1;
  wire [0:0] wire_52;
  wire [0:0] wire_52_0;
  wire [0:0] wire_52_1;
  assign wire_52 = wire_52_0|wire_52_1;
  wire [0:0] wire_53;
  wire [0:0] wire_53_0;
  wire [0:0] wire_53_1;
  assign wire_53 = wire_53_0|wire_53_1;
  wire [0:0] wire_54;
  wire [0:0] wire_54_0;
  wire [0:0] wire_54_1;
  assign wire_54 = wire_54_0|wire_54_1;
  wire [7:0] wire_55;
  wire [7:0] wire_56;
  wire [0:0] wire_57;
  wire [0:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_59_0;
  wire [0:0] wire_59_1;
  assign wire_59 = wire_59_0|wire_59_1;
  wire [0:0] wire_60;
  wire [7:0] wire_61;
  wire [0:0] wire_62;
  wire [0:0] wire_62_0;
  wire [0:0] wire_62_1;
  assign wire_62 = wire_62_0|wire_62_1;
  assign arch_input_enable = wire_62;
  wire [0:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [7:0] wire_66;
  wire [0:0] wire_67;
  wire [0:0] wire_68;
  wire [7:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_70_0;
  wire [0:0] wire_70_1;
  assign wire_70 = wire_70_0|wire_70_1;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [0:0] wire_73;
  wire [7:0] wire_74;

endmodule
