module MUXzm8i (clk, rst, \0 , \1 , \2 , \3 , \4 , \5 , \6 , \7 , Selector, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] \0 ;
  input  wire [7:0] \1 ;
  input  wire [7:0] \2 ;
  input  wire [7:0] \3 ;
  input  wire [7:0] \4 ;
  input  wire [7:0] \5 ;
  input  wire [7:0] \6 ;
  input  wire [7:0] \7 ;
  input  wire [7:0] Selector;
  output  wire [7:0] Output;

  TC_Decoder3 # (.UUID(64'd1969048836624943678 ^ UUID)) Decoder3_0 (.dis(1'd0), .sel0(wire_18), .sel1(wire_2), .sel2(wire_6), .out0(wire_20), .out1(wire_13), .out2(wire_15), .out3(wire_19), .out4(wire_12), .out5(wire_1), .out6(wire_5), .out7(wire_17));
  TC_Splitter8 # (.UUID(64'd1861387493510513996 ^ UUID)) Splitter8_1 (.in(wire_14), .out0(wire_18), .out1(wire_2), .out2(wire_6), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Switch # (.UUID(64'd4405675252321471448 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_2 (.en(wire_20), .in(wire_0), .out(wire_3_7));
  TC_Switch # (.UUID(64'd2626601727990729237 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_3 (.en(wire_12), .in(wire_7), .out(wire_3_6));
  TC_Switch # (.UUID(64'd1330337826708257526 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_4 (.en(wire_1), .in(wire_11), .out(wire_3_4));
  TC_Switch # (.UUID(64'd764843388776523872 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_5 (.en(wire_5), .in(wire_8), .out(wire_3_2));
  TC_Switch # (.UUID(64'd3752377706505052511 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_6 (.en(wire_17), .in(wire_10), .out(wire_3_0));
  TC_Switch # (.UUID(64'd1750255450023985824 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_7 (.en(wire_19), .in(wire_16), .out(wire_3_1));
  TC_Switch # (.UUID(64'd2819839412399577864 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_8 (.en(wire_15), .in(wire_9), .out(wire_3_3));
  TC_Switch # (.UUID(64'd3577968039719068292 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_9 (.en(wire_13), .in(wire_4), .out(wire_3_5));

  wire [7:0] wire_0;
  assign wire_0 = \0 ;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  wire [7:0] wire_3;
  wire [7:0] wire_3_0;
  wire [7:0] wire_3_1;
  wire [7:0] wire_3_2;
  wire [7:0] wire_3_3;
  wire [7:0] wire_3_4;
  wire [7:0] wire_3_5;
  wire [7:0] wire_3_6;
  wire [7:0] wire_3_7;
  assign wire_3 = wire_3_0|wire_3_1|wire_3_2|wire_3_3|wire_3_4|wire_3_5|wire_3_6|wire_3_7;
  assign Output = wire_3;
  wire [7:0] wire_4;
  assign wire_4 = \1 ;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [7:0] wire_7;
  assign wire_7 = \4 ;
  wire [7:0] wire_8;
  assign wire_8 = \6 ;
  wire [7:0] wire_9;
  assign wire_9 = \2 ;
  wire [7:0] wire_10;
  assign wire_10 = \7 ;
  wire [7:0] wire_11;
  assign wire_11 = \5 ;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [7:0] wire_14;
  assign wire_14 = Selector;
  wire [0:0] wire_15;
  wire [7:0] wire_16;
  assign wire_16 = \3 ;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;

endmodule
