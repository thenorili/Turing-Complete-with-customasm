module MUXzm8zp (clk, rst, \0 , \1 , \2 , \3 , \4 , \5 , \6 , \7 , Selector, Disable, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] \0 ;
  input  wire [7:0] \1 ;
  input  wire [7:0] \2 ;
  input  wire [7:0] \3 ;
  input  wire [7:0] \4 ;
  input  wire [7:0] \5 ;
  input  wire [7:0] \6 ;
  input  wire [7:0] \7 ;
  input  wire [7:0] Selector;
  input  wire [0:0] Disable;
  output  wire [7:0] Output;

  TC_Decoder3 # (.UUID(64'd1969048836624943678 ^ UUID)) Decoder3_0 (.dis(1'd0), .sel0(wire_22), .sel1(wire_20), .sel2(wire_21), .out0(wire_3), .out1(wire_19), .out2(wire_13), .out3(wire_0), .out4(wire_10), .out5(wire_9), .out6(wire_7), .out7(wire_5));
  TC_Splitter8 # (.UUID(64'd1861387493510513996 ^ UUID)) Splitter8_1 (.in(wire_11), .out0(wire_22), .out1(wire_20), .out2(wire_21), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Switch # (.UUID(64'd4405675252321471448 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_2 (.en(wire_3), .in(wire_16), .out(wire_4_2));
  TC_Switch # (.UUID(64'd2626601727990729237 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_3 (.en(wire_10), .in(wire_1), .out(wire_4_7));
  TC_Switch # (.UUID(64'd1330337826708257526 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_4 (.en(wire_9), .in(wire_14), .out(wire_4_6));
  TC_Switch # (.UUID(64'd764843388776523872 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_5 (.en(wire_7), .in(wire_17), .out(wire_4_5));
  TC_Switch # (.UUID(64'd3752377706505052511 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_6 (.en(wire_5), .in(wire_6), .out(wire_4_4));
  TC_Switch # (.UUID(64'd1750255450023985824 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_7 (.en(wire_0), .in(wire_2), .out(wire_4_3));
  TC_Switch # (.UUID(64'd2819839412399577864 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_8 (.en(wire_13), .in(wire_15), .out(wire_4_0));
  TC_Switch # (.UUID(64'd3577968039719068292 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_9 (.en(wire_19), .in(wire_12), .out(wire_4_1));
  TC_Switch # (.UUID(64'd3191703730251323901 ^ UUID), .BIT_WIDTH(64'd8)) Output8z_10 (.en(wire_18), .in(wire_4), .out(Output));
  TC_Not # (.UUID(64'd3697959477816005703 ^ UUID), .BIT_WIDTH(64'd1)) Not_11 (.in(wire_8), .out(wire_18));

  wire [0:0] wire_0;
  wire [7:0] wire_1;
  assign wire_1 = \4 ;
  wire [7:0] wire_2;
  assign wire_2 = \3 ;
  wire [0:0] wire_3;
  wire [7:0] wire_4;
  wire [7:0] wire_4_0;
  wire [7:0] wire_4_1;
  wire [7:0] wire_4_2;
  wire [7:0] wire_4_3;
  wire [7:0] wire_4_4;
  wire [7:0] wire_4_5;
  wire [7:0] wire_4_6;
  wire [7:0] wire_4_7;
  assign wire_4 = wire_4_0|wire_4_1|wire_4_2|wire_4_3|wire_4_4|wire_4_5|wire_4_6|wire_4_7;
  wire [0:0] wire_5;
  wire [7:0] wire_6;
  assign wire_6 = \7 ;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  assign wire_8 = Disable;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [7:0] wire_11;
  assign wire_11 = Selector;
  wire [7:0] wire_12;
  assign wire_12 = \1 ;
  wire [0:0] wire_13;
  wire [7:0] wire_14;
  assign wire_14 = \5 ;
  wire [7:0] wire_15;
  assign wire_15 = \2 ;
  wire [7:0] wire_16;
  assign wire_16 = \0 ;
  wire [7:0] wire_17;
  assign wire_17 = \6 ;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;

endmodule
